Description:    Concept of classes data type with example 
************************************************************************/
//ADD_CODE: Declare a class called "simple" with properties i and j of int data type
//          and write a task called printf to display the properties i and j of the class

  
program simple_class;
 initial
   begin
    //ADD_CODE: Declare two handles to the class simple as obj_1 and obj_2
    
    //ADD_CODE: Create object for the handles obj_1 and obj_2
    
    //ADD_CODE: Access property i using obj_1 and initialize it to 2 and 
    //          Access property i using obj_2 and initialize it to 4
    
    
    //ADD_CODE: Call the task printf using obj_1 and obj_2    
    
   end
endprogram

