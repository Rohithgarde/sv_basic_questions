module packed_and_unpacked();

// ADD_CODE:declare a packed array packed_array of 8 bits and initialize it to 8'hAA

// ADD_CODE:declare an unpacked array unpacked_array of 8 bits and initialize it to '{0,0,0,0,0,0,0,1}


initial 
 begin
  //ADD_CODE:display the 0th element of the packed array
  
  //ADD_CODE:display the 0th element of the unpacked array
  
  //ADD_CODE:display the whole packed array. Is it possible???
  
  //ADD_CODE:display the whole unpacked array. Is it possible??? 
  
  #1 $finish;
end

endmodule
