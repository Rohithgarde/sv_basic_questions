
Description:    Concept of class inheritance and constructor with example 
************************************************************************/
//ADD_CODE: Write a class called base with property "value" of type int 
//          explicitly override the class constructor - function new() in the class base 
//          and initialize the variable value to 3 inside the function new()




//ADD_CODE: Write a class called ext which is extended from class base with property "x" of type int 
//          explicitly override the class constructor - function new() in the class ext 
//          and initialize the variable "x" to 5 inside the function new()



    
program constructor1;
  initial
   begin
//ADD_CODE: Declare and create object for handle "e" of the class "ext"
   

//ADD_CODE: Display the variables "value" and "x" using the object "e"
    

   end
endprogram
