module associative_array ();

// ADD_CODE:Declare an associative array as_mem of type int and index type int

// ADD_CODE:Declare a local variable i of type int for manupilation


initial begin
  // ADD_CODE:Add element to the associative array as follows:
  // in the 100th location store value 101
  // in the first location store value 100
  // in the 50th location store value 99
  // in the 256th location store value 77



  // ADD_CODE:Display the size of the associative array
  
  // ADD_CODE:Check if index 2 exists
  
  // ADD_CODE:Check if index 100 exists
  
  // ADD_CODE: Display the value stored in first index
 
  // ADD_CODE:Display the value stored in last index
  
  // ADD_CODE:Delete the first index
  
  
  // ADD_CODE:Display the value stored in first index
 
  #1 $finish;
end

endmodule
