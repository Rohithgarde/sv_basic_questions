module dynamic_array();

// ADD_CODE:Declare a dynamic array mem of 8 bits


initial begin
  // ADD_CODE:Allocate the dynamic array for 4 locations
  $display ("Setting array size to 4");
 
  // ADD_CODE:Initialize the array with 0,1,2,3 values
  $display("Initialize the array with 0,1,2,3 values");
  
  // ADD_CODE:Doubling the size of dynamic array, with old content still valid
  
  // ADD_CODE:Display the current size of the dynamic array
  
  // ADD_CODE:Display the each value and the location of the dynamic array
  
  // ADD_CODE:Delete all the elements in the dynamic array
  
  // ADD_CODE:Display the current size of the dynamic array
  
  #1 $finish;
end

endmodule
