
Description:    Concept of shallow copy with example 
************************************************************************/

program shallow_copy();

//ADD_CODE: Write a class "A" with property "j" of type int and initialize it to 5



//ADD_CODE: Write a class "B" with properties "i" of type int and initialize it to 1
//          and declare handle "a" for class "A" and create object for it
 



initial 
  begin
//ADD_CODE: Declare a handle "b1" for class "B" and Create an object for it
  

//ADD_CODE: Declare a handle "b2" for class "B" 
  

//ADD_CODE: Make a shallow copy of "b1" to "b2" 
   

//ADD_CODE: Display "b1.i, b2.i, b1.a.j, b2.a.j"
  

//ADD_CODE: Now change the value of "i" in "b2" to 10
  

//ADD_CODE: Display "b1.i, b2.i, b1.a.j, b2.a.j"
  

//ADD_CODE: Now change the value of "j" in "b2.a" to 50
  


//ADD_CODE: Display "b1.i, b2.i, b1.a.j, b2.a.j"
  

  end
	
endprogram
	


